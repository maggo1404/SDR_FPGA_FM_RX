--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.09 Education"
--Wed Mar 01 19:18:13 2023

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.09_Education/IDE/ipcore/FIFO_HS/data/fifo_hs.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.09_Education/IDE/ipcore/FIFO_HS/data/fifo_hs_top.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
OAPgg63lQSwlr3ye+vA1rsf1rQ8jEHWY1r9gUsJNuAGPRJL8R4EJzv3ODHGEkyCZDWPGUuuKR1nr
NlvQYi+h8IBf0FuzqbIlXAj5gbg1yNixwvx6X2J3CcH/Yyc8sJRA/G3VfQANc4Pc8J5QTMBhuFDk
FVBVQu/EhlnJYH2x9T75BpHBDNgxVKxijtL3UevtdGHZ/HGUJWy9KAqx6ESun+jUntCe+yZeKKrm
wYGH3EDyQwvR/Fw1ikRmnnfp+ZdO9e/HaVkXEAxS728Hgp3FqbuzA6WBi7MYr3qV1Ct21iva1OOp
2/RJNzRrxrUgwdMw0PDhB8zEau8DDHH70nJyAg==

`protect encoding=(enctype="base64", line_length=76, bytes=12000)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
5uQDz6VioPZxdzMGKtix7TAECgUqf9qQ49NhYZCiEae0aahYQjEBMwvdUC0gG7CsxUEMY7z2g1ay
XFoG/bajveeL0oihL63XOeiIWhAGcmmRBB+p+Z4r5Jeez5sZNCn2LEMjLMtDBb6/Hw/XoFl+AQiC
8v28IZSraSgeCG6RPT9gCAEvMc3EdsFf/3j4S9EDcIdnNJMtOv5VtCZe4mTBMOmXhV1oGFL2Vmmv
vKX+frxx3LLkx/1KnXNNWahBFJwfuVtCDtu79AqCiLKXULnZ8yvxs2WyhLxoXc56Ok1wi8WG8XJ4
g41UAj3F4/OAWshFMroiFF4oXD6m/AUJMQYuCuEv7iOSB73nNe2WTYO6GVHfU79b3Bjt8fqMx3AF
b7D3PIk4HMvz8HKPGtOq5LMdKzQiLFENfo3iGqxyhc92qESSPqdz+A13G4XAO9AHYe+vCinNqiSf
EydIUc6SHd7c56v0m5RtBWM2QxgCq69hKDDQeQHFHBUaTUMRVEJaOofhOSLog7DgxpixeDcigdAx
UYp3GQ7o7mRVo6Vm4cNqzMZFit62kypQZ6xYtBIHREWEqeU6QePvuij7a0lmf40skDLLXsDAE5Xi
svvJQ8+chx/7qqSE1dnXxg3ZgQkwTrtSurWQVqCZDW0RVbBDB/Tw+pLvq0P4Ktbq76ruGnaAQ87X
nuIzqr1L2QyXJZr6YyEB1HPYOzFq+6Jm1CGxMxRWBZAkGozxm+yQovtzSUehfZehe5Srz0rK5Tbz
TQp07Zo7KWfRxQwxnEnCfleN/CHte8JkYrp3D0rVZ6SXdmC9j/z9z+twUtPCSRZUVgVU+F94H4gm
qzfzbg9qqlroWxl4w5POoc3rIOb0Zmv/Hefq+IxlmXLUK1bNn5knXj27U0lVV2t/2S0cfb5xOy7N
/RL/wghxPNGWiupgY/MUThnAXT6oqbv58Nw9cs10OptItBp/zcI04czxwyHGjVZROZCtIeVNyKC9
av4ClXkZon3PLSdr8LLWdDuihn0Z6ZlDaHpKdR4/8TYsh59soS+rPFlxWp9Z8/XXOpx8sP6MyLo1
OkRZ5gwpSd4qf9NuI+xGEm3hR2Os7kpBfc4O8DNP2EoM94RKYg9MOKhkhh2cFx95W3dCxyJ+qB/e
ALBOAUlZPM75WO426Ppb8N3FAEtEJot0MPwx6/21hhDF22WwmtGNE2dbgb34JjD7dsb5h4s1MECR
HHWA2zQrVu46rfpKjWJJrOcyTSNK9sP+8uUhKElOk81Kehz10qy+oEpb/y5ZV5FQsnBou8fEbAwE
PkaBTQbDubNIcRwl5b8GgAuyiXEiEXYNeQcd5dJM2Gl+81o51ah6AaW4gjRXBIo6vtPdToIAJ8B9
cDwCTGZwyFU+mr85DR6p8LgebqbdCj8ZH1dUN00+m2VMJEkgbaRmmeyT/c8vshkLkqxvcBOhZJ25
SXwhGE9/P/6c2YPPD+USVhUUM5ROfWun3ZsXQ6a8b4AfHB7j3LHClWC7soGqEOjfQh4We5385lVf
4qQGo2wloEBHK00yZwI+2bp9puDPvHPUlDznLJ7C1ByEONxJB06miXN73taVmoCrvwrHOrSJ0MNI
6yX06hcO5WY7I9oZv13R9j6NzXYEXdsEbk8fVy+iJh4fdQW2DAzNlRGtfpeET6xUFFbc2dT1vD6v
7hX4Jkn+3ZIb6t59fwrlK/MA59tg21XfflzcieRoQLIej7DR+Hrf2DBDMMkrCxbtIo5B/ON3S6j2
RgrFFj/x3Ql23bLVqEYwaLrGj2DEI0SYDAjQ0Ej2pMpd+odDvRdbCw7kMas7R/W+GxiEBRUl3dVL
Twid0Q9ZSFw2q9ZaZtE8pgKGOAQBC0Zc9HXHNrDS9zTO8JLkxyXJ7+dRcztN9S36wt9MGNY5A9WM
grWgZDtv6I4lQlbCAnSlXRzRDCGJCZqvYBxJlFjPSlQrJmkwPUuXr95JLKPgbGmgbQlvZsdYGrCT
Szxnfn6bx4hgDSVs8km2jD1jL4XYei8T+HR1qgzXbXroM4Mlb7NpQ3vanlFANMPQdh1fpbEQOOpa
mIaSBML3KDLBEtP2t1VYSnj2L7y+XhLji2nBMQCY6p+4q1GR9bUL2riDHQPV4kZf7VAWubc6C+Lx
Xa8m/HWuIqIqcmSmp1ZLqBYi6qnRuQU5aC0v3yLgs7LYtvWTLjdcvfn6/XE/ia9jgs9ydv4cf0hD
pgtTBu9Rmy0IQ4m3QD/F2UbaMzSxBLFRVWqwnP9Etw4U9tUmU63OScB8Tu5jVhcUtvS4SW+nGFyx
WM4MRoSd5uSyZ0x4KbooPgcUqH3/+UKoCGruBbji7Dx8pZPbzE7kPARySDVXCG5Nc0mm2c6D3U9U
Rn02owWYcSSDUZYSPGb/svZVcQPPNShT46E2yDro9518DsAS4IDqyV0nSRCPXFZRTtgr6zZzGiOK
XgqG2ix4pExER4kAowfvWCDmy23cZDbIINq4OtMx3tetmTwVicCxdbxdfR1QBvEaE0KUQ6qEfQo3
glTJt8HN/EoQjKYd7dIBg2YktJ0BM4cvmXZmIWTLnlmOVgD8ejZuEiZvSlyEqEv0xgpIzr9PGQ4j
y9pGSp3RKnjZXCrK8K3bdNGCkQaL35pO7WtBJEVnNHzzWy3aWuhUHlw/RTR6E9Dp3fTmmusxR6Ic
JWsrcsaaQer5770j2WAmIQyzcuvFIov2wGHAtlbP+++buj2uAUU+P+TE/Yb0JlFWquyj856HUvTz
S9IqhExY2t2J7zZgL0NAu/xiZk1IhPG1Xe8lZrse1xTgGi+Txei6yhop8AMp5/0nMYU91fbbQe8g
mXg5gWGzCx7W0Sz4v/tCR81ojk/ZPsl5GPxL4gAR0CLrGKBMt2gunO0VUfNcn/85ndNXIhyOWzzk
6LUJQ5NDV+hHvcYVnlgEU4qBb5toXs1pOmF6zZDjbNG1ua7TnmNMxyESUVNkGnj8IGRPg1aVx4Sz
nfcFlrZLRgwjhEOt6ahohsRs9K+uTy/wMh82QAv7k/rGxqsFzUULWfKx2fxNJDdKYcnGWsWJM9ko
DBFh5dDHZiqeG6I1EQRDIApubSoNc2kr/95OOtbSSsBUsgMS2FzNFfwd9Ka/JLoJ6jsOAHy3/SRo
d7L2dROb0vjSmN2472Kb1kbCZsWQveJEIQBsfNg+orwX6urwIndYCsQaKAquOJR58/YHd1eHV2ek
zegJoZrFHo3VJVRVhfRaPyOS4b96aS2DkHAIBoMS4x92Co8v0CtVSXJgsfkysV2itLNHLnseaY0u
cCtwNp0sEW8PL7WByIvNWIGrZOrtGgb6BHV0AvCVOseUXmqedJJWqb/Oz8I129+86SiCMg6E3s2h
07+SlhD2UBzbzxEH+8FOiciuRloCU720cCzafMZALiKk5x88RPKwbrleSjuMfTPL0P5aWuB2kbDj
ePdzR/Z3jsZUL7RVk/vs9+Jw+s6nik7GK6zZ++LY8Xju93PXdT+nXL921sIlRXw04y4FXTEe5w79
9WY00yZebD1OinMBPq2f0Cm100ILsjOQ75RUXSTzBREqEFbt6vboVjB/fKiPTb5lBoRMzzfIHslV
MZFdNY/shbe5dePbUc5k99gzYmYRXr0TFykL8GQCv+NnweWj/XRqlmI7FE6vzDY08E4kHQ0YoT4R
+U3JrwIvuwz7Vzq5+uon74TLGop3ChbM/hDYWbkap6ONaouJIDOjCr/oE14Rvn5cl4o0+RAwSuCJ
Ke/A1c0SwqJXJ37+DIDKctupAn9b6yuM3SHOpc3GZcezAr/2nOvImZN/OjTy/AWfVwZ7S8eAogzo
m+SlQSIjUVwUlTdZDNwn8X1342wE+UHy/e6WtuGf3UYPTn/EHnO8rwS2ASQAjsYpSy31sqrmUHcb
DVEEouhlWyw/myMQJy78fGvr42kIRa2C6JL9waVqzp+J73mwR6Nm6bpr7jKkt8Dga8YmtCg9CGAf
FetkW/2bP8VahktcVukSg9zNQFc0EaqJ8dk8xXH9fWDAvvb4+LGO2tMTdX/N7LUcNw34m6VWznfv
w1pB8gAUqwuGDDbHmBh/6sZI4I4LC+Ud2E4P4VMuQ54lKHdExOImJ8DO09hPnwMXO1tJq9GWYKbE
PLtxHYoHgwi0zVaiaarLvZEwoasJ6dCypTflLIIfQD3FtRFnT3/qsJ3ehYer0eUl7uN74eEqYT6o
7YGRDKxHv6tf9up93kZodEjmh251XRPOlsgIBKNjvshKxbe20umMidnIVFbs+YTCNDCiIQx7sJON
8+DOHZRrbT+FmjzcHo3NyQCJfq6L2bxwIf9sVh+NJHD9ZhBqejogJY9BlbLTboK3JeFFYhnSY60v
PddVtY3kvH4F5aqRuvDI+qwk2vP5bK3jVECl6ugq8BVWDNhWPJDndfY+pVZTI9W8u6n9YHKM30N0
IGQcgmZKUYjIhYWK8+Wpeh5y24V2IWKcUKXBToELF+Q/JunPVnxY49A0gb7K9CddYq1V9N/xoFCB
NZMqtof1YAuOXoGetGUY8d1kXeqKXgbbZk6vMkLQsq6EjxkLKlPN2GwF4eentviFqccLlQadZiZw
rqj3AMnIcBhPZTn+Yo1PvQctv6SAXxW3GL/fDoW/2uIkWhS/vgZdI6vJqV7Ja1hZAkYyNO0sDBUN
hhocw9lSB1M367QkIDYjPFRbyK2cQQqhXRxJ40U5+8XsH9BYU7X/jc8k/doS/8kBADr4pDaWyWiK
GBr+ajJPjobn9mV0WNX2oa7me9scjNgOc3eBW7/J3J55N8nDrWVMop9q3nFsLyowfWThjg+2wzjH
P5zc5pRWHpOqCz1jtypjkqymtNfoc1AgJc/OGT2qs1Q0cLxE3+SX3ovLj/XdOtMg5MEpX7WxovL7
+n3g2LjSQsAuGuCHb5VwvR6utM8rKIai82qnQSRUNeLcBxGVyueMCLgANKAmCJESyIkQ/a9ArKxx
fDtOiP7uyPRSeZYwwjW0sTesoTNpRn8AZZkN/+sb2smnd08NJieY3AfTTYwjqT2oS9SppF1Xd5yL
q0pJSKDPvclYPGma74z6fi7KtAOvIxjKaThO3do/vgE4V26cYMh5OK64GmibbYLnFdVPcJZSpN9D
bV+151Q89IPLoqs5AoIA/IDybyuJPD26hlE821m5Zi2gTijJrJ1jda+FRf1H0iR6M8BMz8ge34Tl
5b2G7RbN8FtbVqvglEljJ/080YG4aL053N5991W/l4tgH1RbkGydbrljzD0HyUpyBu0IB6dZ/Ium
G4OtIxW6IwpU2EtC9KIEu4I4jtxyCU6fdhpEh7btEtaQmo2ysLcVhRhLzD/03yMCDkaiVFxGE4vn
YduFlBYL6vxgfqNmkqeX0EXeSx7AcbIWSoIenuPIefxZHlKC+05BAKb3AteQux+73l9oIHH6rF2Y
JidjXHNmrX8W8CRkD/tUIxLNYKdJtNyfUXaCGAYizQmI3oZEtkOg5zv5zWnapGMLiho/VRSvr4Vr
rdGrBeTa96fpUJy6xwILzLqPHQubb8bE3O93wF9t8Slht7BhgK2pz5tkZ8LB53bY1YlccvrY6Og/
/L+cCfxAQmwLGmbPOggT9qt6aIcwknU0uvbsESTDLGZrbZUbZx0Q/RV+XfDzdvTL5Ra+bw7ce15Y
2n87g7NPjkwsnCE54q8B1WSlV+A2gOfqC0agQc9vJ6Eg6xY1CzyyRuTv0LXF8g3uQcfxHrYk/vti
NnODZOevpw/dUueskzNxg63nxEDaMzfw4h0d0Fqjfu+sfSv+A4supdwaayFmFtRIvbx8TkGHcYkr
Y5Ef4fmgg3PChj9BwKyZsxXa/EKcjsoIcljscSlvhJBq4fPEYy9uB+w+cODxyMehO2PMM3vG0cPt
Ve6/RHRt6cZZ+SQt0EyMDB6AZLWSdHwykPnCdMhmZT0jdKWPg+YrDCLVPSyjzlgaxLnhsDqRLfVk
ppPVd0WOh2BNk2DyVBaZkdQV6II8G72mZREErMy6WTj2RPHPeYySDlnjDM3XFCq9Wetr1JfyFL61
6UoEx0g4HOxlhwqeAxn97U53nLGWce1jo5vqPhl5bssOHFf/kBi5wRleO9D0MZoPyLh6AeHUrhT9
xSId+FIPJqYMkbABfHOTb5X8HTIs5hRlV803QQYS4M3bIdC343MkjDDH50WEweidavJ1bl3UWGnW
rTF9vxF8egj+IwhwR3If6jq+sDLQHvRIIGd+Bbm56ELfrRBh+vD1hOqHY3yLvUa4scS80oy93L7A
q32IsgshtQPORg57ycBew5TweEQQlIxGBOy6ikO17mr62tqkn/FSyNig0TJJirDXg96MQ5aGWtvt
WZY/yvV+jZTg10QFqKbEV/2uPcPbFKyfsWJWkrT9MmJ6CsOsgykAtYJ8VISckTLR9JCgdtkksGTX
0VfXKcj7cufCj/3EhOxVFEVyhFlzpOzSAI/2235dDjzr9ntyXqRYBGmGs0eBjQvo1E94+H9yR+3K
7aEICDHY5b1V0KPACzxoeHWNbCBZWG7Mfgfs81NDGYwO+i+jV8r4xSdFrUBQ/k1KlPprq9RJ0Het
1na66frH6YuzoS0iPNUHPe6hhzY+AY2I9tLvf/ebchriji0Ms0UCx1kpg/Xbynmsup52ZM4GhGeW
twb8EIU8S2gUnYDCMxmAVTwJd467CVwZNP9aa1CpvF3XC2kR1Hp5IhNQsk3k1A1sfxm2XuREJnH7
hoGsRkfCutTkYOk5LZUSNUJSjfNmlq+Kykw/5G/IdWg2S7kV8JMJoc1VnQZdLo+Qx+oShIrmbqRu
6dJkbtYV7d7V0kJ2WEafNIkHO9TqgtTg85y35yCDJEbE7m7cWkVPWhtI0KQvRAXnu50DZtnNlSpg
WZXjyd24CILTReQhH2uPREaPAkbqMxsfHOLeRLLyeuuVo7qqaoFbSYYHnfGjZfMUBZOgZsdji580
vdig8URmEfL00Dvg7LHfVO7aW0GYOdLhPNNVvnSp1Js/blU2kQ5nEJEJe3XL4NYoq2QN7SYhN6ws
SgjnfS/qcudkbRIzZHcMJumv5nJDy7/6AABe8jL1E6LIXzXVTZjb7OIWTSNa1Zp8AfKQxXKpt7kZ
4NXBP1UoKoTcrmO7siFaXgGT09A9klbD5sKTcBI68cMHbpDXdtafzFeseEFLtkiUMybF4/pt6OiZ
F1P9VWY9frpgDjqqpTgietfcS4Bj6ebnC+A87RGQ6ac9ivCXW9k2MtxIbkLAYtHWwhLv9LmnEnz6
YtVUvhbaGutVk6pYdjBONUCPTaM3eJ3XGInBXeoMsKqKLZ1ojZBwggoObLlO6IVlRmPSiOjHoRW9
9wjk3t8KXHMP7/KaXT82aoKL78F2vgwxVlBLXfdI21q/SoqpKmeVTDSm4xC1Lh303QLXCoZ5I1pZ
yojEGO+TS5xwEYdt8sVJohXRGnvd8l9JCsjCyHrvf/N9HFLPIZJCGmXMdF5SNvbViwF6MWw259BR
iNEx1Om98gQy92wwifddDm3NVdDLJUWCBPimY4cpVEA5jJGw+f/Cm4zMqx0IL3ptmeDidjlKC3u+
grDcMbY3FDlvR98/HrYvKDdbUnJENAVFney2DQleSJs/lMsAae5KVcJ7RiioQgu6M/h9jjmAQzrT
xVgeQikjUbfEYOn+ije+3MNcBTbtrTy6863ymcQca+ZheMlGrp4JF785qAMP9CKQszzLa33MHBob
ybnk7wKCfFsi+4fE03yEgbg+X3mFtWQ2ZEaTki6ilc1hin39uzWSLPVN0txAOwuRlVWnTP1WZCO1
EGzMyvc8Fivk0Ed1/DbGdkDQHQe/S1b8c5pzuPeOpbFDH8eCh6xC9yVRWme1aiXIY7kmU0c13EXN
qq9f+g7g9Y81ROFZ7cGSiO7oTCvLoKHqpbIDG6pNVzn9m7ZAb9E60EiKdb9gqIX15rTjTnI75Gqk
1ZNdyL5tWsh3QgSXtdUQC6/iAtW8fI5KAQRE313glfb1z2KemgHMvEJEZDxPyZgHLyep9E4xbbGJ
idvLxizOFC2RNOEMvCFAqGJhtW5m4EGw4cdqDxAEe5t1bM6gNnm1aAHpEXT79tvLfunzJMWRmBs4
awDU9JSc9o8ri+e2oZYRpyIF82tQTBx9cLUNhgoTh7cItxW9p/7FRgaC3629+4CL/2DnltazcpZV
+EC0iV8IKjDq4iwuLXZ+FqDcRoSD3hUe5skzqT0XljiNX/lriQ6TD4E3ZnBfyFEM7GWJUHRVlvKW
1G3oB5hCgOnoq4leEtA2nZnqEtOMP7IzmgzY2RhIUoL5RiUI6o27crf5esx0NxFRmvUPRL0b/2/k
gOn0ZjTPKGV1d2hjNJImupnIKUAadt5sKXwMsJ0fNzqdO+x0kBxIfmxrn/9JQ3z7YdNMjafj1kMH
Bhvj1mVJHEe9Vm/MWzerOnj/yD599jx+Hkbm7ZIHijS8Ng5ql7jozSyNztyApF8ScVxMWPxq1jQH
7RLJXlIUbVilcvrhizCNW71uQucni3iJsIsiitZ7osIBCP8P5Vv0PWtkwBEJCgoqzSggllzeVsgI
EUHXlm9a264wTMVIz6TViHdljzbMM0nBH0JFpiB/TFnWKWW4AMCsNkaoEAnkKYmN8QhQi+Alll86
L+k9IqDk7qLc6z0SAanb6kYOmQufRhPUakNCqvs5KZ/jTns1eyMwoGE4P4F06P12KnZGQuCdTKZD
YWchDGUv97REPpH4KuLKjxKWQ1QqMp6NEUw+BV0FQmVqoSDqppqbLtkdvBMWY2+4Cz3Jk/ASUaDd
DuTolvh7hkp1aaHGuRpfKRTaKAblPDkFndLsDVAqRLBr3crfTQE85RIRKlkrSvUc1wZsgZW/zcuv
U6sMG8cy0lXfpD2LqxerPtjk+UD5/0E6IJ4U2uQjAQ41ALVvAFIoiPAXb1ywIs6XkWkmw2RU4qdD
CqXAW+LC8cAoYftcYnzp3k6g9yyRE3/E8gIBSJ5MgC7CNyS6r8dXj8v6+wMD8KDwZcHOvQOzDqac
0dOSfK7njH4vW4VeYITBPKPuBAXFUxW1thjYMG0dHGrUQxjG0lEi+zQqlKPhQxJVipwiRDdy9B2H
vJTniRT0tq7Lvzk9z353eNFIDhP5wZmSFdKhEh2y1tIeOu24IXAErLCn5ZE3u7In0TmQcqH3iHnV
0cZE4hPtSWI19LwHmOfyu/p18k0Xu7Zs/wue7y73dyLypw6Sqx/Ltu/IAP6ZofPBDy79u0WNOqq4
SKMtU5LyS8YsSC1M5ajWbE10PJ5VmdhjPu/ZUJEwPP8twZUGtNkbikTFwFncjmc/Qf2udjPDCKMh
k1vMnhAY2Mcm4wGSkcPvb68TKsGgzEGOZ2ClahBWz4L6yOHUzQhXMBY3HS5Pwe/XV7ao2DChDP5k
/OkZgu+QtS3phn8jk0H3L+f8V9w9Mf/FiSk2JHK1YJL3B/uR/329vPmE3jGYn+agQ3Wv7XGzOYkA
runE1YPmw7e4RtL3xdziLktRvMxjkmR6ysq7cd0uZsq5AWQMa2J+5+LqoilNJi1yq8bZNjGoiHH7
Qzy7Wc8WPCSRUG8nR8wi5+SGlm6mDDRSLudv8e4lkoiVyt5pO2GddupxAT1LbqktS+WYWFr2YgVm
xXVTnATKgHpqyOr12nYP15BRkmUwaH9n/YXChCrva/1R1pv3fv9yaIn772mC0mVE6YL6UaZIugv0
4Rn9XdPyxjZmwG6f8bfXipBxokju4YtfHMExSjWZHwtc7zzv3yjzcxw5V++GPo3MWQFJunVpFlLG
8bxQ2HyM/u8lnNcXfZlmmIo9eGZDViWJJSQDll9Cb5ziTtudlY7XlPcN4UaAhtM+IWqE7hoO1rot
+8OOxLY3J5lv11O4voC8iNX1VUhsOkM+yg3YfMZPYfcGT+5WuH9oz3aSC7s6f6bkblImqkI4RZeJ
EYHGWxUJT/F0S08di6/EM3KJMcQGPkluj1IrgyKuM7apdaZYy3qFab/f5mTlRLJBefYVgr+AwvK3
HDyaHL9aL8/9ujMWjCyLYA9sHW/MWPPuPM6AiBjcorm6psMbwBC+HBlE1efm0oxkEgMwJeAWQFCe
9TvWIrJK5iKzGp7amonPskUrH5TTaII2BQq2aXX0p+3utBw5o2b/vc6FzxdAtdVLiQlwyUZKuU4h
ML+1zZbuFeF387iwJptgmHTo4nGDqlt/MH/5Yhh5TCTr6WzC/8EERVKPCJM0IuHm6ocISeQRnxSG
OuObu2eC8XGvyUL2q60vApk2lX06nRoRoAZnJLIS6yNDCRnsUxNvvxiLBqk7jZhTvcxrTdebnkGW
0G9+VatLeFm2muhK9i8fEqY+5R7IPt3kydA2vG9BIdzIcORGjDxDJDEJ+dzz5xnqAFotfIKtnaGf
Sl94CzVJy9FFPxbDq+V5db2vXGfIvT0QgrUgcQg30hRLxmLkSD41EiXiYycv4NcMfwFS0dtRYJZX
FzluhTzg+lEp5QD65mI+Q8jhDR6hO24ySiSAOQodGCOUDP0ECSXRwg/tdx1pI/WA5Px9k5pMauvW
ZtbVn93su/Sqv69aEsNCx0CEC0/0KJyei8mrv5i+ZVpgLRWkGRmVncMdhMsEz4sQ3b2mTw0963oc
VMY61lyJuV79DgVFtmoY4scCIr5IlrBavwTw93yx3RbE1/j5hL2qAj1zGFGJEfoOWl2+gZ4rTOV2
5/WzZ++U8oguXJsJ/OV7mR2VLASdDXcdYoNb/oGGEUI7gSRorxs+Fg6HcAMHolsYN/yyyIzrmH3i
1HddGBSGyW0IQml/6ksPMfP22ZysEtIHA8Da4uOCpamDgWY936Bs2JZugeQx1rPhTS3Ix5PdSa6M
pKGL9ZOSsbPonEfMRZ2oAsry7aRvCsUb+614qk+/bcX7hYSSBmXz+gH8PCuGfAEQWONUIFx7yH2C
qrK/PyU51Rqh5IMKzjhpvKKZ9qeug0TwvhBQRH+BLTeFt+dGApT1qBpQlVI1sZ/hj116ihZkVo0U
tJTtehcvVFcIlFHH/5cV7WI5PCY5X1TkbqYU2tZyqaPjlh4GlLp0HK116FIcpnpD4ykaZACbqrVo
Lw8xIDBSSSuHNNfiLlXsaPgDJNCKJLpJS543sDnpi5gt66cd0u3FprwX0oyG/rHcF6N6aqB1QMfm
RWNfusSFUrgFVCsmQByFwXJMiMEqBywYoFsq/ierMBLfCzyB4de5x/FxjogIG1wIpuAvIIstoCG5
akOM7Ws3aTl5D0BU5tzqzctV+F0U6i12Z2RgYVnbnaJuB9njQCiNAGvL4DRm+gZU3JTUCZ/S2p3I
aJSVRdJBOOMb9RympkB71KmBm0SCeoEFXaZckXj4Qj1Q9G1/LHGGSKK+ejItQZ2ckExX9fADgS0J
UlAlTDESOlFYVIdtapMZViu1+2tu4t2zuggirytanKzCclB3Cyu9d06SXGYapwAG5CinIHmu9+q7
qmhd+s7gecuQHe9bEtBjkbeP/SYzWrrOmH9NTj6DyH9STrMd6GKemLOaQ+KEegZWqx1GnLJqYHiv
QUDvB6PilRlLjuhIJW4CPO/k4gNZRpird0niM2X9im5bCiK5YCeBmveIBcaFuEl1CzgjzJmm1brF
pbI957pOtcCLh77IpaexooY6Q8Wdr8Xuht99UNbHzHRqcFFtw/G05VkYMlbfHFp75ytmqzkOgcrr
ByJWE8x0+NWuxnNT7DmyzsELBHPWnTTeiynX2TfokalgIg8Bf7I6sSrGYt2YWdzcFlz1IjtC9eTm
WDR66qVpPRPStsuchuP4s0VRBov1mL/3Rs58u5ChWWZWlw0bKl07PtnB7TiBhRNcETquEBJv0jRq
27svzaM+w7NtRgNl4EQ/6o6fsqDOPu7qknu/0c3GLTKt+ZDeuFbaaiqvKUqM4p7A8AXJPVYOp36E
yDdqrJ3ZlPcAYDPql5ygi1KYDWb7cQdkmc1TVsZXkLSKH2ilHEpiGS/W5Wc7Bj+QocEkYEfDCt2e
DFTkaHbJVBJ1LGZ7QQS3/zf15H6gZ7Sy4zSmdTAisNad1/Tod/xwhDd1rqTw3gBeD9DyFIJuOesA
lXTPQDaDhdvMmJksfc69sTXsPjI3SA8Qjw7UCfXsKQxV0Q7O8qNbXgsGLJ3myHOu9G2gTVNkZBVt
m2/92dZQEtYYDoaGTUkWNxovdRVDlNZmr5L7RTLFVb49gt/FpHdayK1jTd0PnQB0MyvwkDVXaBUy
5nX1PAZBUabMUU11paF5bTDpnjzDu1zj4uJ2WzTHfO3OwdnbWpsSSDKwkPtS3LP4XvtHaK6umrs2
DCIktwx/0gjbkNhJIasXKIZLX5pNKEJ1KFhRZANS7P5uvtJpdnP2ec/myKptfM1R9PqFZozwO6/Z
A+EY5R9u31rg9SrqlFXykJTfCoI6ullfcQLTtqq7WYxErPN7QSAJGhdIloWiJok3DE/vq6pgqhqb
ekioTCYgZDbOsY76sONdcj6eUKZaLr0mUyRMteq1QLkby3mVJsI99TaG1wbNL9+saPfu6Gu0lF9C
7R8NMK/5CZ3j0k+nPVeYFxkxmxV3m+bfXftFHb0NoxPvdy6bN7WktuvXyFvR38ZuN/92MVEcFNyf
UOQ52aignsEW77q3DB2GpFafBdgG9U+1jjkjzQlPiO/T9vJ/2oVBg5RA7/VgmUamRz4Tx4/nXVTy
x8Q9bQ/tV9fAQRVu1u4li26ekLFYN00qiErOSE2iu+9ARmo1uvMY0WQ/uaP1r9D+0oAqHk7o92n5
CG8OR3E7aGLbiZM9GMapaJC6xAstZ8EC1lwCgwdmDQyAOhT0UrL0MIsMxFdo/BfCVMPAJOhWQHHi
O3oqcanANWjkcLTqgHOTiNNIDR48y4IF6b0DfPwZsEYnBRHYNdDhLIjzR2UD+2tuzsBB7YnM3sS1
ZXdORj9ZFW35KyGJmKpwYPFhsVKU8/egOZE/cpyxGK3Qt2leUH7r3LoGOiYl63IOW6PuNNg/EIRZ
3Izsq89vOreM8zbRW9jl3Vk0ZKGuN0zIQGZgYA05hUR0Gon4adR/PhodzOehDwQ3N8TRIg0VbyGC
LXlLm9h9dIcY9Y69IrNhn9EL4tVqcT5ymm2/zBILRdxx57u0vo+jOyjjg/iMtrvESlwgSwiB+RRP
vYiUh4ipBWXFJ3eDLMWNqI4CfkbIFG4cBYpNMyFqIiOTLDKoYE7JQ4FEFHhkFxvbn0cNdPnognw5
4z+9zaQ2IVVIJ1XE2Q5nluLNx/Cs+HMAcAamceIYANH2zbz5pGJGIaJbWgIyqPRZieMu3yQyqnY6
wDE/iXJUyj6azzkuDmlyoh3xgs23epHDoK1mNAa6SH9xWluGO5Vjx4SltIxICEv5mvCLwQLekzoJ
RbF4rz3+fJUgOmLkMHz15XxmQmyl9GKeO7wHqvE2XpMFcqf0O4zQOzr/1WBgoXN01jUJZaikGlWt
fNEObbxM3o0bvmjdYpc7scTg1MBaKBDvZj9COEU4JpuCIa8ru/johjolOnRl5jbaPvznJbWduIjQ
14n88tGgyFt3VhPv6IJkhj5I+wJ7jf0YZ+t0DikMXdRFrj9+AbqKMmL7ZlX1OsvOU06dx/T4PfnT
ZujtrQFEAy5ue97B0KpZ/0k3yT4MIzsf+QNjJHqnREZ9AVOZNQb8JO4ifFZY6NkNyBI9xfeBM/yD
zDjqvEi4cP9hCA61gJUalmmRvNokciLAlln2r4L6iy6sP5ohSXAI95oqRAr/NDuI2bLov96zaXCe
6UPhV50Boeusgp8ySKWZKoPDGWFIsKSu/Z0eYpuWSri+b2W1sNZNSdNyeukrMPsxSO7AxWZijqfM
9ZGOZpuW5zeukgi4x4E4GeUhk7BWlzP4yiI4gCMvz6XhWFqNuVPYBolexQdkAJ+gat85VwiCET/0
bFu6KRIEzc46pXWcZoo9PeJqOl/vIpApZGKyF3kJhvjWsgqh1sPDJAJcHy2/7KFbhzPwlVWb470D
vniryMmyStw3CkBkrqW92tTzjbZyqbn0uKbGuXUdU+vEHAbhVMed8YlZG9y9DeRgDCzIWyQXiX0S
sYLoTy/bYJ3a0711kBlrwtLxZvKBDt7iENGqUxg8YK8U/h+dh3oqwjCiR8Y5VGKZGA0E5riZlppQ
hSrKAQ153k8VH/c/+e+XVXqILIQ8tZz2W6eTXjM453JBZMikCaeVScY5lqH4cP75hh2zL+GunDLs
WsOLdDo0MfPJyDE/bYMfGWCW4/HCOk2AlQWq9nlLgdTFL3nJ8fSlKJGiXCU6qI9/Xq2t6WJQatgc
AekOZP8+OR8nMVebMYsOiH6RDdq1twcRBh1IMPWz6QULNlg5rCrpbdzj6LX4wARioLSBsHj5mYMd
wWn9hRP9T0Anfx1ahU9JfuvZaakpe6zrcaFayN3fpnND1I9P3CqU0+06qk2oUOP1TwXNyj5Rqdmy
qQG7OtC7OFC1KLSrnc5Fum4Fw0Kxv63F6cAf1s6xq8DHQWqkHpH9lx0G1Sjh+uRTQQ3wJG4YRFjh
fM/ZGIWak4aTjxMe/avGotr7mTn6zxaZ0uEVdtfQx3PTE5uz4T0LbvGhcavK7XSCgcAofcLLjCft
yGPtbBzw/snRFtq7lw51Pca683VVxxSvJ5fSZiZVQpXUf+EunDX/Uk8b/wNDwaqto7Vy5OtWiAWK
NmtlnUpAvlOQII/KXuFWzie2cZrfQtNL40J0rJnRZpFItBngsIZbqZo/lN3MGZEhPaaQOY1QFcds
CqpFHAECzwAL+dHlpi2cw7kw691jrx8qPdC3WLmKwi+bAMVNf/uG915dkM+Xt1kKE9Xf05Y7mkke
dx97T+LZs2UBiB3IT4jHNDWWAGGfkfrDpZt4tMTO9OiwTbKPfbOxR9L28qcCNzghC2CN+ylJSe+k
YI69jFdnR0ArGudlJski5zbiKerjH6/oO69A/504fiUmf2M1qQQV6it0wg+SSiQ40YkmzGEi0DUa
AftF2zidlhieOozHRQlrIzn1zvSE4GNvOsJ9IRLkBfyIK3WVpTUjftsJBwjRT7JLuJqh5y8I7cfs
HpK0KC0vG3Qtb/ee/03s3lTelA8SlPrpAtrG2qlpUB5J1S6L/l+TvbqGz+7S6R+y6FizsfFirsjw
Tv8vGVM9Oi8okRZlHfnmzn1fbIBNTBhp6ZFYgYeEK00HRMOeXzCYtIn0VJ6nGjuB8f5g3uuZf0Xk
0ypXFsNqiIqCwhJD3DUygJAHaj90+tGgzSq0trruMddQFGhJfWOlQTfAQHnh2CVtGD7FEwca1M/2
F2bPZDm93OYUTx0Y7QLI+YcecfZCDjb5D206ypxdfC2ndR7dJQXpFWrPJNNMRm+xmP5AXOCFQHSq
ViT8CeqLU/YJL8FjfZlD3Bi65PCWsaYPrnM2Iv0f2E2h9Qn9LTVK9lH3WaQ8iTyE8Fz7WNUAXzWO
oIsLrrU+rG7MtqCVMGvUtxcev8CRhWfnfTygyNSzpS7AHciyMIBinT74agkLEM+oFunoHX4s3B4H
xu1jN8OFFtrPyJJYaFLf/7N8bT7ZTaKd1qV21Ynd29pyTncGlIB/QWWIKXGxrvpiz/3CBMnbkDh0
C0tDqZdvMJRS1ByrL+vVvv7hVnez59fzl2wFulITItiofOlYHwUmpWuy74TmoHnpaif5VhqAPRi4
Nmltu+/kbsGcjDqoItahs0M8PygIZiEUcKfX16rXQmGRry0C0a1IkbzAvNlk5e9/pJDBqLVRCCGW
Pc+4OoDyQQBl7NXCVwFLUKzAr90Gh6z7HayeZLeHUxQD1QfT/1C1OxrvV3DavhXRXu2/Huyt2wXI
ZM4pvKkvWNDWVKvWD3CaLU1s8G2UfATlXFB8J0AHqqHJxeAmI1/aoqH770qr3ETljFsUyXwmQ7ma
tkRColAhHmR7NQMOpowfAp3Ue24MLZG9RjyuxOapDSUaB/xSKtI8h+Xy18Tr+5xuz1CZ/7Y+781R
644KnsdT7W9at2b6P4B9xqnqmgyegKX8fvTwFjvirvKLwVGo6L9PGyfrFPBy19j4Le7QCmUn32vI
gfaztX3obIsasowU/ZV6Uwxb2ymZ89Lxu0CHe7lA
`protect end_protected
